library verilog;
use verilog.vl_types.all;
entity SignExtend_vlg_vec_tst is
end SignExtend_vlg_vec_tst;
