library verilog;
use verilog.vl_types.all;
entity mux8_1_testbench is
end mux8_1_testbench;
