library verilog;
use verilog.vl_types.all;
entity mux32x32_32_testbench is
end mux32x32_32_testbench;
