library verilog;
use verilog.vl_types.all;
entity mux32_1_testbench is
end mux32_1_testbench;
