library verilog;
use verilog.vl_types.all;
entity decoder3_8_testbench is
end decoder3_8_testbench;
