library verilog;
use verilog.vl_types.all;
entity comparator32_vlg_vec_tst is
end comparator32_vlg_vec_tst;
