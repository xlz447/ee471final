library verilog;
use verilog.vl_types.all;
entity decoder2_4_testbench is
end decoder2_4_testbench;
