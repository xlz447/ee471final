library verilog;
use verilog.vl_types.all;
entity comparator6_vlg_vec_tst is
end comparator6_vlg_vec_tst;
