library verilog;
use verilog.vl_types.all;
entity decoder5_32_testbench is
end decoder5_32_testbench;
