library verilog;
use verilog.vl_types.all;
entity mux2x6_vlg_vec_tst is
end mux2x6_vlg_vec_tst;
