library verilog;
use verilog.vl_types.all;
entity c_tb is
end c_tb;
